-- Elementos de Sistemas
-- by Luciano Soares
-- Register32.vhd

Library ieee;
use ieee.std_logic_1164.all;

entity Register32 is
	port(
		clock:   in STD_LOGIC;
		input:   in STD_LOGIC_VECTOR(31 downto 0);
		load:    in STD_LOGIC;
		output: out STD_LOGIC_VECTOR(31 downto 0)
	);
end entity;

architecture arch of Register32 is
  -- Aqui declaramos sinais (fios auxiliares)
  -- e componentes (outros módulos) que serao
  -- utilizados nesse modulo.
component Register16 is
port(
		clock:   in STD_LOGIC;
		input:   in STD_LOGIC_VECTOR(15 downto 0);
		load:    in STD_LOGIC;
		output: out STD_LOGIC_VECTOR(15 downto 0)
	);
end component;

signal signal1, signal2 : STD_LOGIC_VECTOR(15 downto 0);

begin
	bite1: Register16 port map(
		clock  => clock,
		input  => input(15 downto 0),
		load   => load,
		output => signal1);

	bite2: Register16 port map(
		clock    => clock,
		input => input(31 downto 16),
		load => load,
		output => signal2);		

	output <= signal2 & signal1;
	
end architecture;