library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Or16 is
	port ( 
			a:   in  STD_LOGIC_VECTOR(15 downto 0);
			b:   in  STD_LOGIC_VECTOR(15 downto 0);
			q:   out STD_LOGIC_VECTOR(15 downto 0));
end entity;

architecture arch of Or16 is
begin
<<<<<<< HEAD
--<<<<<<< HEAD
--q <= a or b;
--=======
-->>>>>>> upstream/master
=======

q <= a or b;
>>>>>>> master

end architecture;
