-- Elementos de Sistemas
-- by Luciano Soares
-- Register8.vhd

Library ieee;
use ieee.std_logic_1164.all;

entity Register8 is
	port(
		clock:   in STD_LOGIC;
		input:   in STD_LOGIC_VECTOR(7 downto 0);
		load:    in STD_LOGIC;
		output: out STD_LOGIC_VECTOR(7 downto 0)
	);
end entity;

architecture arch of Register8 is
  -- Aqui declaramos sinais (fios auxiliares)
  -- e componentes (outros módulos) que serao
  -- utilizados nesse modulo.
 component BinaryDigit is
	port(
		clock: in STD_LOGIC;
		input:   in STD_LOGIC;
		load:    in STD_LOGIC;
		output: out STD_LOGIC
	);
	end component;
	
begin
	u1: BinaryDigit port map(clock,input(0),load,output(0));
	u2: BinaryDigit port map(clock,input(1),load,output(1));
	u3: BinaryDigit port map(clock,input(2),load,output(2));
	u4: BinaryDigit port map(clock,input(3),load,output(3));
	u5: BinaryDigit port map(clock,input(4),load,output(4));
	u6: BinaryDigit port map(clock,input(5),load,output(5));
	u7: BinaryDigit port map(clock,input(6),load,output(6));
	u8: BinaryDigit port map(clock,input(7),load,output(7));

end architecture;
-- Elementos de Sistemas
-- by Luciano Soares
-- Register32.vhd

Library ieee;
use ieee.std_logic_1164.all;

entity Register32 is
	port(
		clock:   in STD_LOGIC;
		input:   in STD_LOGIC_VECTOR(31 downto 0);
		load:    in STD_LOGIC;
		output: out STD_LOGIC_VECTOR(31 downto 0)
	);
end entity;

architecture arch of Register32 is
  -- Aqui declaramos sinais (fios auxiliares)
  -- e componentes (outros módulos) que serao
  -- utilizados nesse modulo.
component Register16 is
port(
		clock:   in STD_LOGIC;
		input:   in STD_LOGIC_VECTOR(15 downto 0);
		load:    in STD_LOGIC;
		output: out STD_LOGIC_VECTOR(15 downto 0)
	);
end component;

signal signal1, signal2 : STD_LOGIC_VECTOR(15 downto 0);

begin
	bite1: Register16 port map(
		clock  => clock,
		input  => input(15 downto 0),
		load   => load,
		output => signal1);

	bite2: Register16 port map(
		clock    => clock,
		input => input(31 downto 16),
		load => load,
		output => signal2);		

	output <= signal2 & signal1;
	
end architecture;